// Lab 2
// Created by David Tran
// Last Modified 01-22-2014

//Verilog HDL for "es210",

module flip_me (A,B);

  input A;
  output B;

  not G1(B,A);

endmodule
